//dataflow
module not_gate(output Y,input A);
assign Y=~A;
endmodule
