//gate level
module and_gate(output Y,input A,input B);
and(Y,A,B);
endmodule
