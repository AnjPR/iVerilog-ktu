include "program1.v"
module program1_tb()
reg A,B;

