//gate level
module nor_gate(output Y,input A,input B);
nor(Y,A,B);
endmodule
