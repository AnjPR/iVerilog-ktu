//dataflow
module and_gate(output Y,input A,input B);
assign Y=A&B;
endmodule
