//gate level
module not_gate(output Y,input A);
not(Y,A);
endmodule
