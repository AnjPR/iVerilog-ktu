//gate level
module or_gate(output Y,input A,input B);
or(Y,A,B);
endmodule
