//gate level
module and_gate(output Y,input A,input B);
or(Y,A,B);
endmodule
