//dataflow
module nor_gate(output Y,input A,input B);
assign Y=~(A|B);
endmodule
