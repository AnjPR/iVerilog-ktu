//gate level
module nand_gate(output Y,input A,input B);
nand(Y,A,B);
endmodule
